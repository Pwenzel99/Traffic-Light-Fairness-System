module seven_seg_decoder(o,x);
	input [3:0] x;
	output [6:0] o;
	reg [6:0] o;
	
	always @(x[3] or x[2] or x[1] or x[0])
	begin
		case({x[3],x[2],x[1],x[0]})
			4'b0000: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0000001;
			4'b0001: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b1001111;
			4'b0010: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0010010;
			4'b0011: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0000110;
			4'b0100: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b1001100;
			4'b0101: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0100100;
			4'b0110: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0100000;
			4'b0111: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0001111;
			4'b1000: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0000000;
			4'b1001: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0000100;
			4'b1010: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0001000;
			4'b1011: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b1100000;
			4'b1100: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0110001;
			4'b1101: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b1000010;
			4'b1110: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0110000;
			4'b1111: {o[0],o[1],o[2],o[3],o[4],o[5],o[6]} = 7'b0111000;
		endcase
	end
endmodule
